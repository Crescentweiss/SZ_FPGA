module SZHDPredictor(
  input         clock,
  input         reset,
  input  [31:0] io_in_0, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_1, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_2, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_3, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_4, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_5, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_6, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_7, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_8, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_9, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_10, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_11, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_12, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_13, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_14, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_15, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [31:0] io_in_16, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [4:0]  io_startindex, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [4:0]  io_midindex, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  input  [4:0]  io_endindex, // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
  output [31:0] io_prediction // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 8:16]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] datareconstruction_0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_1; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_2; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_3; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_4; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_5; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_6; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_7; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_8; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_9; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_10; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_11; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_12; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_13; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_14; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_15; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  reg [31:0] datareconstruction_16; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
  wire [4:0] dataprediction_size = io_endindex - io_startindex; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 25:44]
  wire [4:0] dataprediction_left = io_midindex - io_startindex; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 26:44]
  wire [4:0] dataprediction_right = io_endindex - io_midindex; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 27:43]
  wire [31:0] _GEN_1 = 5'h1 == io_startindex ? $signed(datareconstruction_1) : $signed(datareconstruction_0); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_2 = 5'h2 == io_startindex ? $signed(datareconstruction_2) : $signed(_GEN_1); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_3 = 5'h3 == io_startindex ? $signed(datareconstruction_3) : $signed(_GEN_2); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_4 = 5'h4 == io_startindex ? $signed(datareconstruction_4) : $signed(_GEN_3); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_5 = 5'h5 == io_startindex ? $signed(datareconstruction_5) : $signed(_GEN_4); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_6 = 5'h6 == io_startindex ? $signed(datareconstruction_6) : $signed(_GEN_5); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_7 = 5'h7 == io_startindex ? $signed(datareconstruction_7) : $signed(_GEN_6); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_8 = 5'h8 == io_startindex ? $signed(datareconstruction_8) : $signed(_GEN_7); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_9 = 5'h9 == io_startindex ? $signed(datareconstruction_9) : $signed(_GEN_8); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_10 = 5'ha == io_startindex ? $signed(datareconstruction_10) : $signed(_GEN_9); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_11 = 5'hb == io_startindex ? $signed(datareconstruction_11) : $signed(_GEN_10); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_12 = 5'hc == io_startindex ? $signed(datareconstruction_12) : $signed(_GEN_11); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_13 = 5'hd == io_startindex ? $signed(datareconstruction_13) : $signed(_GEN_12); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_14 = 5'he == io_startindex ? $signed(datareconstruction_14) : $signed(_GEN_13); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_15 = 5'hf == io_startindex ? $signed(datareconstruction_15) : $signed(_GEN_14); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [31:0] _GEN_16 = 5'h10 == io_startindex ? $signed(datareconstruction_16) : $signed(_GEN_15); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{59,59}]
  wire [36:0] _dataprediction_prediction_T = $signed(_GEN_16) * $signed(dataprediction_right); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:59]
  wire [31:0] _GEN_18 = 5'h1 == io_endindex ? $signed(datareconstruction_1) : $signed(datareconstruction_0); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_19 = 5'h2 == io_endindex ? $signed(datareconstruction_2) : $signed(_GEN_18); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_20 = 5'h3 == io_endindex ? $signed(datareconstruction_3) : $signed(_GEN_19); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_21 = 5'h4 == io_endindex ? $signed(datareconstruction_4) : $signed(_GEN_20); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_22 = 5'h5 == io_endindex ? $signed(datareconstruction_5) : $signed(_GEN_21); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_23 = 5'h6 == io_endindex ? $signed(datareconstruction_6) : $signed(_GEN_22); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_24 = 5'h7 == io_endindex ? $signed(datareconstruction_7) : $signed(_GEN_23); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_25 = 5'h8 == io_endindex ? $signed(datareconstruction_8) : $signed(_GEN_24); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_26 = 5'h9 == io_endindex ? $signed(datareconstruction_9) : $signed(_GEN_25); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_27 = 5'ha == io_endindex ? $signed(datareconstruction_10) : $signed(_GEN_26); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_28 = 5'hb == io_endindex ? $signed(datareconstruction_11) : $signed(_GEN_27); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_29 = 5'hc == io_endindex ? $signed(datareconstruction_12) : $signed(_GEN_28); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_30 = 5'hd == io_endindex ? $signed(datareconstruction_13) : $signed(_GEN_29); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_31 = 5'he == io_endindex ? $signed(datareconstruction_14) : $signed(_GEN_30); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_32 = 5'hf == io_endindex ? $signed(datareconstruction_15) : $signed(_GEN_31); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [31:0] _GEN_33 = 5'h10 == io_endindex ? $signed(datareconstruction_16) : $signed(_GEN_32); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:{98,98}]
  wire [36:0] _dataprediction_prediction_T_1 = $signed(_GEN_33) * $signed(dataprediction_left); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:98]
  wire [36:0] _dataprediction_prediction_T_4 = $signed(_dataprediction_prediction_T) + $signed(
    _dataprediction_prediction_T_1); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:67]
  wire [37:0] _dataprediction_prediction_T_5 = $signed(_dataprediction_prediction_T_4) / $signed(dataprediction_size); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 35:106]
  wire [37:0] _GEN_34 = io_midindex == io_endindex ? $signed({{6{datareconstruction_0[31]}},datareconstruction_0}) :
    $signed(_dataprediction_prediction_T_5); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 32:43 33:24 35:24]
  wire [37:0] _GEN_35 = io_midindex == io_startindex ? $signed(38'sh0) : $signed(_GEN_34); // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 30:39 31:24]
  assign io_prediction = _GEN_35[31:0]; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 29:30]
  always @(posedge clock) begin
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_0 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_0 <= io_in_0; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_1 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_1 <= io_in_1; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_2 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_2 <= io_in_2; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_3 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_3 <= io_in_3; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_4 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_4 <= io_in_4; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_5 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_5 <= io_in_5; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_6 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_6 <= io_in_6; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_7 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_7 <= io_in_7; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_8 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_8 <= io_in_8; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_9 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_9 <= io_in_9; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_10 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_10 <= io_in_10; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_11 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_11 <= io_in_11; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_12 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_12 <= io_in_12; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_13 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_13 <= io_in_13; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_14 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_14 <= io_in_14; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_15 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_15 <= io_in_15; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
    if (reset) begin // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
      datareconstruction_16 <= 32'sh0; // @[\\src\\main\\scala\\example\\SZ_HD_1parameter.scala 21:35]
    end else begin
      datareconstruction_16 <= io_in_16; // @[\\src\\main\\scala\\example\\SZ_HD_2predictor.scala 17:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  datareconstruction_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  datareconstruction_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  datareconstruction_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  datareconstruction_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  datareconstruction_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  datareconstruction_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  datareconstruction_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  datareconstruction_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  datareconstruction_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  datareconstruction_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  datareconstruction_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  datareconstruction_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  datareconstruction_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  datareconstruction_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  datareconstruction_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  datareconstruction_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  datareconstruction_16 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
